library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity processador_tb is
end entity processador_tb;

architecture rtl of processador_tb is
    [signals]
begin

    [concurrent statements]

end architecture rtl;